library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package polynomial_cfg is
    constant a :positive :=3;
    constant b :positive :=2;
    constant c :positive :=9;
    constant d :positive :=1;
    constant in_bits :positive :=6;
    constant out_bits :positive :=24;
end package polynomial_cfg;
